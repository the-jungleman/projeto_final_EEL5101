library ieee;
use ieee.std_logic_1164.all; 

entity alpha0_mux is port(
    
    alpha_a: in std_logic_vector(7  downto 0);
    end_game, end_sequence, end_round: in std_logic;
    R1, E1, E2, E3, E4, E5, E6: out std_logic);

end alpha0_mux;

architecture arc_alpha0_mux of alpha0_mux is


end arc_alpha0_mux;               
